netcdf input4 {
dimensions:
	y = 5 ;
	x = 8 ;
variables:
	double t ;
		t:units = "days since 2018-12-01" ;
		t:standard_name = "time" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 t = -10 ;

group: group1 {
  dimensions:
  	lat = 5 ;
  	bounds2 = 2 ;
  	lon = 8 ;
  variables:
  	double lat_bnds(lat, bounds2) ;
  	double lat(lat) ;
  		lat:units = "degrees_north" ;
  		lat:standard_name = "latitude" ;
  		lat:bounds = "/group1/lat_bnds" ;
  	double lon_bnds(lon, bounds2) ;
  	double lon(lon) ;
  		lon:units = "degrees_east" ;
  		lon:standard_name = "longitude" ;
  		lon:bounds = "/group1/lon_bnds" ;
  	double time ;
  		time:units = "days since 2018-12-01" ;
  		time:standard_name = "time" ;
  	double q(lat, lon) ;
  		q:project = "research" ;
  		q:standard_name = "specific_humidity" ;
  		q:units = "1" ;
  		q:coordinates = "/group1/time" ;
  		q:cell_methods = "area: mean any_valid_name: mean time: mean bounds2: mean" ;
  	double q2(lat, lon) ;
  		q2:project = "research" ;
  		q2:standard_name = "specific_humidity2" ;
  		q2:units = "1" ;
  		q2:cell_methods = "area: mean any_valid_name: mean time: mean bounds2: mean" ;
  	double q3(lat, lon) ;
  		q3:project = "research" ;
  		q3:standard_name = "specific_humidity3" ;
  		q3:units = "1" ;
  		q3:coordinates = "/group1/time lon_bnds" ;
  		q3:cell_methods = "area: mean any_valid_name: mean time: mean lon_bnds: mean" ;
  	double y(y) ;
  		y:units = "degrees_north" ;
  		y:standard_name = "latitude" ;
  	double x(x) ;
  		x:units = "degrees_east" ;
  		x:standard_name = "longitude" ;
  	double tas(y, x) ;
  		tas:project = "research" ;
  		tas:standard_name = "specific_humidity" ;
  		tas:units = "1" ;
  		tas:coordinates = "t" ;
  		tas:cell_methods = "y: x: mean (interval: 1 degree comment: comment 1 here) t: maximum (comment 2 here)" ;
  data:

   lat_bnds =
  -90, -60,
  -60, -30,
  -30, 30,
  30, 60,
  60, 90 ;

   lat = -75, -45, 0, 45, 75 ;

   lon_bnds =
  0, 45,
  45, 90,
  90, 135,
  135, 180,
  180, 225,
  225, 270,
  270, 315,
  315, 360 ;

   lon = 22.5, 67.5, 112.5, 157.5, 202.5, 247.5, 292.5, 337.5 ;

   time = 31 ;

   q =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;

   q2 =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;

   q3 =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;

   y = 2, 2, 2, 2, 2 ;

   x = 1, 1, 1, 1, 1, 1, 1, 1 ;

   tas =
  0.007, 0.034, 0.003, 0.014, 0.018, 0.037, 0.024, 0.029,
  0.023, 0.036, 0.045, 0.062, 0.046, 0.073, 0.006, 0.066,
  0.11, 0.131, 0.124, 0.146, 0.087, 0.103, 0.057, 0.011,
  0.029, 0.059, 0.039, 0.07, 0.058, 0.072, 0.009, 0.017,
  0.006, 0.036, 0.019, 0.035, 0.018, 0.037, 0.034, 0.013 ;
  } // group group1
}
