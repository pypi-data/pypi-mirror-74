netcdf input2 {
group: group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890 {
group: group67890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890 {
    		:attr_short_2345678901234567890123456789012345678901 = "This attribute name would be flattened as 255 character long." ;
    		:attr_exact_23456789012345678901234567890123456789012 = "This attribute name would be flattened as 256 character long." ;
  		:attr_long1_234567890123456789012345678901234567890123 = "This attribute name would be flattened as 257 character long." ;
  		:attr_long2_234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012 = "This attribute name would be flattened as 416 character long, and with hashing the path would be 255 characters long." ;
                :attr_long3_23456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234567890123456789012345678901234 = "This attribute name would be flattened as 417 characters long, and with hashing the path would be 256 characters long." ;
    }
  }
}
